`timescale 1ns/1ns

module  tb_hdmi_colorbar();



endmodule
