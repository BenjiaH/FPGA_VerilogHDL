module  led
(
    input   wire        key_in,
    output  wire        led_out //无逗号
);

assign led_out = key_in;


endmodule
