module example
(
    input   wire

)