module  
(

);



endmodule
